module Controlador_display_7Segmentos_tb; 
    reg [3:0] i_Datos_0;
    reg [3:0] i_Datos_1;
    reg [3:0] i_Datos_2;
    reg [3:0] i_Datos_3;
    reg i_Reloj;
    reg i_Reset;
    wire [6:0] o_Segmentos;
    wire [3:0] o_Anodo_4_Bits;
    
    controlador_display_7segmentos uut(
     .i_Datos_0(.i_Datos_0),
     .i_Datos_1(.i_Datos_1),
     .i_Datos_2(.i_Datos_2),
     .i_Datos_3(.i_Datos_3),
     .i_Reloj(i_Reloj),
     .i_Reset(i_Reset),
     .o_Segmentos(o_Segmentos),
     .o_Anodo_4_Bits(o_Anodo_4_Bits)
  );
  
initial 
begin 
  i_Reset= 0;
         i_Reloj  = 0;
        i_Datos0= 4'd1;
        i_Datos1= 4'd2;
        i_Datos2= 4'd3;
        i_Datos3= 4'd4;
        #2 
        i_Reloj =1;
        i_Reset = 1;    

        
  end 
        always
       #1 i_Reloj  = ! i_Reloj ; 
endmodule

